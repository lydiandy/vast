module main

import vast

fn main() {
	file:='./demo.v'
	vast.json_file(file)
}