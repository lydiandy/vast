module main

import v.token
import v.parser
import v.table
import v.ast
import v.pref
import os

const (
	version = '0.0.1'
)

fn main() {
	if os.args.len != 2 {
		println('unknown args,Usage:vast demo.v')
		return
	}
	file := os.args[1]
	// file:='./example/demo.v'
	if os.file_ext(file) != '.v' {
		println('the file must be v file')
		return
	}
	if !os.exists(file) {
		println('the v file does not exist')
		return
	}
	apath := abs_path(file)
	json_file(apath)
}

struct Tree {
	root         &C.cJSON // the root of tree
	table        &table.Table
	pref         &pref.Preferences
	global_scope &ast.Scope
}

// generate json file with the same file name
fn json_file(file string) {
	ast_json := json(file)
	json_file := file[0..file.len - 2] + '.json'
	os.write_file(json_file, ast_json)
}

// generate json string
fn json(file string) string {
	t := Tree{
		root: create_object()
		table: table.new_table()
		pref: &pref.Preferences{}
		global_scope: &ast.Scope{
			start_pos: 0
			parent: 0
		}
	}
	ast_file := parser.parse_file(file, t.table, .skip_comments, t.pref, t.global_scope)
	to_object(t.root, 'ast_type', t.string_node('ast.File'))
	to_object(t.root, 'path', t.string_node(ast_file.path))
	to_object(t.root, 'mod', t.mod(ast_file.mod))
	to_object(t.root, 'imports', t.imports(ast_file.imports))
	to_object(t.root, 'scope', t.scope(ast_file.scope))
	to_object(t.root, 'global_scope', t.scope(ast_file.global_scope))
	to_object(t.root, 'stmts', t.stmts(ast_file.stmts))
	// generate the ast string
	s := json_print(t.root)
	return s
}

// basic type node
fn (t Tree) string_node(val string) &C.cJSON {
	return create_string(val)
}

fn (t Tree) number_node(val int) &C.cJSON {
	return create_number(val)
}

fn (t Tree) bool_node(val bool) &C.cJSON {
	if val {
		return create_true()
	} else {
		return create_false()
	}
}

fn (t Tree) null_node() &C.cJSON {
	return create_null()
}

// todo
fn (t Tree) typ_node(typ table.Type) &C.cJSON {
	if typ == 0 {
		return create_string('')
	} else {
		// type_str:=t.table.get_type_symbol(typ)
		type_str := t.table.type_to_str(typ)
		println(type_str)
		return create_string(type_str)
	}
}

// ast.File node
fn (t Tree) mod(mod ast.Module) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Module'))
	to_object(obj, 'name', t.string_node(mod.name))
	to_object(obj, 'path', t.string_node(mod.path))
	to_object(obj, 'expr', t.expr(mod.expr))
	to_object(obj, 'is_skipped', t.bool_node(mod.is_skipped))
	to_object(obj, 'pos', t.position(mod.pos))
	return obj
}

fn (t Tree) imports(imports []ast.Import) &C.cJSON {
	imps := create_array()
	for imp in imports {
		obj := create_object()
		to_object(obj, 'mod', t.string_node(imp.mod))
		to_object(obj, 'alias', t.string_node(imp.alias))
		to_object(obj, 'pos', t.position(imp.pos))
		to_array(imps, obj)
	}
	return imps
}

fn (t Tree) scope(scope ast.Scope) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Scope'))
	to_object(obj, 'parent', t.string_node(ptr_str(scope.parent)))
	children_arr := create_array()
	for s in scope.children {
		mut children_obj := create_object()
		to_object(children_obj, 'parent', t.string_node(ptr_str(s.parent)))
		to_object(children_obj, 'start_pos', t.number_node(s.start_pos))
		to_object(children_obj, 'end_pos', t.number_node(s.end_pos))
		to_array(children_arr, children_obj)
	}
	to_object(obj, 'children', children_arr)
	to_object(obj, 'start_pos', t.number_node(scope.start_pos))
	to_object(obj, 'end_pos', t.number_node(scope.end_pos))
	to_object(obj, 'objects', t.objects(scope.objects))
	return obj
}

fn (t Tree) objects(so map[string]ast.ScopeObject) &C.cJSON {
	obj := create_object()
	for key, val in so {
		to_object(obj, key, t.scope_object(val))
	}
	return obj
}

fn (t Tree) scope_object(node ast.ScopeObject) &C.cJSON {
	obj := create_object()
	match node {
		ast.ConstField { t.const_field(it) }
		ast.GlobalDecl { t.global_decl(it) }
		ast.Var { t.var(it) }
	}
	return obj
}

fn (t Tree) var(it ast.Var) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Var'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'is_mut', t.bool_node(it.is_mut))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'is_used', t.bool_node(it.is_used))
	return obj
}

// stmt node
fn (t Tree) stmts(stmts []ast.Stmt) &C.cJSON {
	stmt_array := create_array()
	for s in stmts {
		to_array(stmt_array, t.stmt(s))
	}
	return stmt_array
}

fn (t Tree) stmt(node ast.Stmt) &C.cJSON {
	match node {
		ast.Module { return t.mod(it) }
		ast.Import { return t.import_(it) }
		ast.Comment { return t.comment(it) }
		ast.ConstDecl { return t.const_decl(it) }
		ast.FnDecl { return t.fn_decl(it) }
		ast.StructDecl { return t.struct_decl(it) }
		ast.EnumDecl { return t.enum_decl(it) }
		ast.InterfaceDecl { return t.interface_decl(it) }
		ast.Attr { return t.attr(it) }
		ast.HashStmt { return t.hash_stmt(it) }
		ast.CompIf { return t.comp_if(it) }
		ast.GlobalDecl { return t.global_decl(it) }
		ast.DeferStmt { return t.defer_stmt(it) }
		ast.TypeDecl { return t.type_decl(it) }
		ast.GotoLabel { return t.goto_label(it) }
		ast.GotoStmt { return t.goto_stmt(it) }
		ast.AssignStmt { return t.assign_stmt(it) }
		ast.Return { return t.return_(it) }
		ast.ForCStmt { return t.for_c_stmt(it) }
		ast.ForStmt { return t.for_stmt(it) }
		ast.ForInStmt { return t.for_in_stmt(it) }
		ast.BranchStmt { return t.branch_stmt(it) }
		ast.AssertStmt { return t.assert_stmt(it) }
		ast.UnsafeStmt { return t.unsafe_stmt(it) }
		ast.ExprStmt { return t.expr_stmt(it) }
		ast.GoStmt { return t.go_stmt(it) }
		ast.Block { return t.block(it) }
		ast.ComptimeCall { return t.comptime_call(it) }
	}
}

fn (t Tree) import_(it ast.Import) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Import'))
	to_object(obj, 'mod', t.string_node(it.mod))
	to_object(obj, 'alias', t.string_node(it.alias))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) position(p token.Position) &C.cJSON {
	obj := create_object()
	to_object(obj, 'line_nr', t.number_node(p.line_nr))
	to_object(obj, 'pos', t.number_node(p.pos))
	return obj
}

fn (t Tree) comment(it ast.Comment) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Comment'))
	to_object(obj, 'text', t.string_node(it.text))
	to_object(obj, 'is_multi', t.bool_node(it.is_multi))
	to_object(obj, 'line_nr', t.number_node(it.line_nr))
	to_object(obj, 'pos', t.position(it.pos))
	// to_object(obj, 'same_line', t.bool_node(it.same_line))
	return obj
}

fn (t Tree) const_decl(it ast.ConstDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ConstDecl'))
	field_arr := create_array()
	for f in it.fields {
		to_array(field_arr, t.const_field(f))
	}
	to_object(obj, 'fields', field_arr)
	to_object(obj, 'is_pub', t.bool_node(it.is_pub))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) const_field(it ast.ConstField) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ConstField'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'is_pub', t.bool_node(it.is_pub))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'comment', t.comment(it.comment))
	return obj
}

fn (t Tree) fn_decl(it ast.FnDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('FnDecl'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'return_type', t.number_node(int(it.return_type)))
	to_object(obj, 'is_deprecated', t.bool_node(it.is_deprecated))
	to_object(obj, 'is_pub', t.bool_node(it.is_pub))
	to_object(obj, 'is_variadic', t.bool_node(it.is_variadic))
	to_object(obj, 'is_anon', t.bool_node(it.is_anon))
	to_object(obj, 'receiver', t.field(it.receiver))
	to_object(obj, 'receiver_pos', t.position(it.receiver_pos))
	to_object(obj, 'is_method', t.bool_node(it.is_method))
	to_object(obj, 'rec_mut', t.bool_node(it.rec_mut))
	to_object(obj, 'language', t.number_node(int(it.language)))
	to_object(obj, 'no_body', t.bool_node(it.no_body))
	to_object(obj, 'is_builtin', t.bool_node(it.is_builtin))
	to_object(obj, 'is_generic', t.bool_node(it.is_generic))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'body_pos', t.position(it.body_pos))
	to_object(obj, 'file', t.string_node(it.file))
	arg_arr := create_array()
	for a in it.args {
		to_array(arg_arr, t.arg(a))
	}
	to_object(obj, 'args', arg_arr)
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	return obj
}

fn (t Tree) anon_fn(it ast.AnonFn) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('AnonFn'))
	to_object(obj, 'decl', t.fn_decl(it.decl))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	return obj
}

fn (t Tree) struct_decl(it ast.StructDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('StructDecl'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'is_pub', t.bool_node(it.is_pub))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'mut_pos', t.number_node(it.mut_pos))
	to_object(obj, 'pub_pos', t.number_node(it.pub_pos))
	to_object(obj, 'pub_mut_pos', t.number_node(it.pub_mut_pos))
	to_object(obj, 'language', t.number_node(int(it.language)))
	to_object(obj, 'is_union', t.bool_node(it.is_union))
	to_object(obj, 'attr', t.string_node(it.attr))
	f_arr := create_array()
	for f in it.fields {
		to_array(f_arr, t.struct_field(f))
	}
	to_object(obj, 'fields', f_arr)
	return obj
}

fn (t Tree) enum_decl(it ast.EnumDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('EnumDecl'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'is_pub', t.bool_node(it.is_pub))
	to_object(obj, 'is_flag', t.bool_node(it.is_flag))
	to_object(obj, 'pos', t.position(it.pos))
	f_arr := create_array()
	for f in it.fields {
		to_array(f_arr, t.enum_field(f))
	}
	to_object(obj, 'fields', f_arr)
	return obj
}

fn (t Tree) enum_field(it ast.EnumField) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('EnumField'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'has_expr', t.bool_node(it.has_expr))
	to_object(obj, 'expr', t.expr(it.expr))
	return obj
}

fn (t Tree) interface_decl(it ast.InterfaceDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('InterfaceDecl'))
	to_object(obj, 'name', t.string_node(it.name))
	str_arr := create_array()
	for s in it.field_names {
		to_array(str_arr, t.string_node(s))
	}
	to_object(obj, 'field_names', str_arr)
	m_arr := create_array()
	for m in it.methods {
		to_array(m_arr, t.fn_decl(m))
	}
	to_object(obj, 'methods', m_arr)
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) attr(it ast.Attr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Attr'))
	to_object(obj, 'name', t.string_node(it.name))
	return obj
}

fn (t Tree) hash_stmt(it ast.HashStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('HashStmt'))
	to_object(obj, 'val', t.string_node(it.val))
	to_object(obj, 'mod', t.string_node(it.mod))
	return obj
}

fn (t Tree) comp_if(it ast.CompIf) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('CompIf'))
	to_object(obj, 'val', t.string_node(it.val))
	to_object(obj, 'is_not', t.bool_node(it.is_not))
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	else_stmt_arr := create_array()
	for s in it.else_stmts {
		to_array(else_stmt_arr, t.stmt(s))
	}
	to_object(else_stmt_arr, 'else_stmts', else_stmt_arr)
	to_object(obj, 'has_else', t.bool_node(it.has_else))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) global_decl(it ast.GlobalDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('GlobalDecl'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'has_expr', t.bool_node(it.has_expr))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) defer_stmt(it ast.DeferStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('DeferStmt'))
	stmt_array := create_array()
	for s in it.stmts {
		to_array(stmt_array, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_array)
	to_object(obj, 'ifdef', t.string_node(it.ifdef))
	return obj
}

fn (t Tree) type_decl(node ast.TypeDecl) &C.cJSON {
	match node {
		ast.AliasTypeDecl { return t.alias_type_decl(it) }
		ast.SumTypeDecl { return t.sum_type_decl(it) }
		ast.FnTypeDecl { return t.fn_type_decl(it) }
	}
}

fn (t Tree) alias_type_decl(it ast.AliasTypeDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('AliasTypeDecl'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'is_pub', t.bool_node(it.is_pub))
	to_object(obj, 'parent_type', t.number_node(int(it.parent_type)))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) sum_type_decl(it ast.SumTypeDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('SumTypeDecl'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'is_pub', t.bool_node(it.is_pub))
	t_arr := create_array()
	for s in it.sub_types {
		to_array(t_arr, t.number_node(int(s)))
	}
	to_object(obj, 'sub_types', t_arr)
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) fn_type_decl(it ast.FnTypeDecl) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('FnTypeDecl'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'is_pub', t.bool_node(it.is_pub))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) struct_field(it ast.StructField) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('StructField'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'comment', t.comment(it.comment))
	to_object(obj, 'default_expr', t.expr(it.default_expr))
	to_object(obj, 'has_default_expr', t.bool_node(it.has_default_expr))
	arr := create_array()
	for a in it.attrs {
		to_array(arr, t.string_node(a))
	}
	to_object(obj, 'attrs', arr)
	to_object(obj, 'is_public', t.bool_node(it.is_public))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	return obj
}

fn (t Tree) field(it ast.Field) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Field'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) arg(it table.Arg) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Arg'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'is_mut', t.bool_node(it.is_mut))
	return obj
}

fn (t Tree) goto_label(it ast.GotoLabel) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('GotoLabel'))
	to_object(obj, 'name', t.string_node(it.name))
	return obj
}

fn (t Tree) goto_stmt(it ast.GotoStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('GotoStmt'))
	to_object(obj, 'name', t.string_node(it.name))
	return obj
}

fn (t Tree) lambda(it ast.Lambda) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Lambda'))
	to_object(obj, 'name', t.string_node(it.name))
	return obj
}

fn (t Tree) assign_stmt(it ast.AssignStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('AssignStmt'))
	i_arr := create_array()
	for i in it.left {
		to_array(i_arr, t.ident(i))
	}
	to_object(obj, 'left', i_arr)
	e_arr := create_array()
	for e in it.right {
		to_array(e_arr, t.expr(e))
	}
	to_object(obj, 'right', e_arr)
	to_object(obj, 'op', t.number_node(int(it.op)))
	to_object(obj, 'pos', t.position(it.pos))
	lt_arr := create_array()
	for s in it.left_types {
		to_array(lt_arr, t.number_node(int(s)))
	}
	to_object(obj, 'left_types', lt_arr)
	rt_arr := create_array()
	for s in it.left_types {
		to_array(rt_arr, t.number_node(int(s)))
	}
	to_object(obj, 'right_types', rt_arr)
	to_object(obj, 'has_cross_var', t.bool_node(it.has_cross_var))
	return obj
}

fn (t Tree) var_decl(it ast.Var) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Var'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'is_mut', t.bool_node(it.is_mut))
	to_object(obj, 'is_arg', t.bool_node(it.is_arg))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'is_used', t.bool_node(it.is_used))
	return obj
}

fn (t Tree) return_(it ast.Return) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Return'))
	e_arr := create_array()
	for e in it.exprs {
		to_array(e_arr, t.expr(e))
	}
	to_object(obj, 'exprs', e_arr)
	to_object(obj, 'pos', t.position(it.pos))
	t_arr := create_array()
	for s in it.types {
		to_array(t_arr, t.number_node(int(s)))
	}
	to_object(obj, 'types', t_arr)
	return obj
}

// fn (t Tree) return_stmt(it ast.ReturnStmt) &C.cJSON {
// obj := create_object()
// to_object(obj, 'ast_type', t.string_node('ReturnStmt'))
// to_object(obj, 'tok_kind', t.number_node(int(it.tok_kind)))
// to_object(obj, 'pos', t.position(it.pos))
// e_arr := create_array()
// for e in it.results {
// to_array(e_arr, t.expr(e))
// }
// to_object(obj, 'results', e_arr)
// return obj
// }
fn (t Tree) for_c_stmt(it ast.ForCStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ForCStmt'))
	to_object(obj, 'init', t.stmt(it.init))
	to_object(obj, 'has_init', t.bool_node(it.has_init))
	to_object(obj, 'cond', t.expr(it.cond))
	to_object(obj, 'has_cond', t.bool_node(it.has_cond))
	to_object(obj, 'inc', t.expr(it.inc))
	to_object(obj, 'has_inc', t.bool_node(it.has_inc))
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) for_stmt(it ast.ForStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ForStmt'))
	to_object(obj, 'cond', t.expr(it.cond))
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'is_inf', t.bool_node(it.is_inf))
	return obj
}

fn (t Tree) for_in_stmt(it ast.ForInStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ForInStmt'))
	to_object(obj, 'key_var', t.string_node(it.key_var))
	to_object(obj, 'val_var', t.string_node(it.val_var))
	to_object(obj, 'cond', t.expr(it.cond))
	to_object(obj, 'is_range', t.bool_node(it.is_range))
	to_object(obj, 'high', t.expr(it.high))
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'key_type', t.number_node(int(it.key_type)))
	to_object(obj, 'val_type', t.number_node(int(it.val_type)))
	to_object(obj, 'cond_type', t.number_node(int(it.cond_type)))
	to_object(obj, 'kind', t.number_node(int(it.kind)))
	return obj
}

fn (t Tree) branch_stmt(it ast.BranchStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('BranchStmt'))
	to_object(obj, 'tok', t.number_node(int(&it.tok)))
	return obj
}

fn (t Tree) assert_stmt(it ast.AssertStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('AssertStmt'))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) unsafe_stmt(it ast.UnsafeStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('UnsafeStmt'))
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	return obj
}

fn (t Tree) go_stmt(it ast.GoStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('GoStmt'))
	to_object(obj, 'call_expr', t.expr(it.call_expr))
	return obj
}

fn (t Tree) block(it ast.Block) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Block'))
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	return obj
}

fn (t Tree) comptime_call(it ast.ComptimeCall) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ComptimeCall'))
	to_object(obj, 'method_name', t.string_node(it.method_name))
	to_object(obj, 'left', t.expr(it.left))
	return obj
}

fn (t Tree) expr_stmt(it ast.ExprStmt) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ExprStmt'))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

// expr
fn (t Tree) expr(e ast.Expr) &C.cJSON {
	match e {
		ast.IntegerLiteral {
			return t.integer_literal(it)
		}
		ast.FloatLiteral {
			return t.float_literal(it)
		}
		ast.StringLiteral {
			return t.string_literal(it)
		}
		ast.CharLiteral {
			return t.char_literal(it)
		}
		ast.BoolLiteral {
			return t.bool_literal(it)
		}
		ast.StringInterLiteral {
			return t.string_inter_literal(it)
		}
		ast.EnumVal {
			return t.enum_val(it)
		}
		ast.Assoc {
			return t.assoc(it)
		}
		ast.CastExpr {
			return t.cast_expr(it)
		}
		ast.AsCast {
			return t.as_cast(it)
		}
		ast.Type {
			return t.type_expr(it)
		}
		ast.SizeOf {
			return t.size_of(it)
		}
		ast.PrefixExpr {
			return t.prefix_expr(it)
		}
		ast.AssignExpr {
			return t.assign_expr(it)
		}
		ast.InfixExpr {
			return t.infix_expr(it)
		}
		ast.IndexExpr {
			return t.index_expr(it)
		}
		ast.PostfixExpr {
			return t.postfix_expr(it)
		}
		ast.SelectorExpr {
			return t.selector_expr(it)
		}
		ast.RangeExpr {
			return t.range_expr(it)
		}
		ast.IfExpr {
			return t.if_expr(it)
		}
		ast.Ident {
			return t.ident(it)
		}
		ast.CallExpr {
			return t.call_expr(it)
		}
		ast.OrExpr {
			return t.or_expr(it)
		}
		ast.StructInit {
			return t.struct_init(it)
		}
		ast.ArrayInit {
			return t.array_init(it)
		}
		ast.MapInit {
			return t.map_init(it)
		}
		ast.None {
			return t.none_expr(it)
		}
		ast.ParExpr {
			return t.par_expr(it)
		}
		ast.IfGuardExpr {
			return t.if_guard_expr(it)
		}
		ast.MatchExpr {
			return t.match_expr(it)
		}
		ast.ConcatExpr {
			return t.concat_expr(it)
		}
		ast.TypeOf {
			return t.type_of(it)
		}
		ast.Likely {
			return t.likely(it)
		}
		else {
			// println('unknown expr')
			return t.null_node()
		}
	}
}

fn (t Tree) integer_literal(it ast.IntegerLiteral) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('IntegerLiteral'))
	to_object(obj, 'val', t.string_node(it.val))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) float_literal(it ast.FloatLiteral) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('FloatLiteral'))
	to_object(obj, 'val', t.string_node(it.val))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) string_literal(it ast.StringLiteral) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('StringLiteral'))
	to_object(obj, 'val', t.string_node(it.val))
	to_object(obj, 'is_raw', t.bool_node(it.is_raw))
	to_object(obj, 'language', t.number_node(int(it.language)))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) char_literal(it ast.CharLiteral) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('CharLiteral'))
	to_object(obj, 'val', t.string_node(it.val))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) bool_literal(it ast.BoolLiteral) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('BoolLiteral'))
	to_object(obj, 'val', t.bool_node(it.val))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) string_inter_literal(it ast.StringInterLiteral) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('StringInterLiteral'))
	v_arr := create_array()
	for v in it.vals {
		to_array(v_arr, t.string_node(v))
	}
	to_object(obj, 'vals', v_arr)
	s_arr := create_array()
	for s in it.expr_fmts {
		to_array(s_arr, t.string_node(s))
	}
	to_object(obj, 'expr_fmts', s_arr)
	e_arr := create_array()
	for e in it.exprs {
		to_array(e_arr, t.expr(e))
	}
	to_object(obj, 'exprs', e_arr)
	et_arr := create_array()
	for e in it.expr_types {
		to_array(et_arr, t.number_node(int(e)))
	}
	to_object(obj, 'expr_types', et_arr)
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) enum_val(it ast.EnumVal) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('EnumVal'))
	to_object(obj, 'enum_name', t.string_node(it.enum_name))
	to_object(obj, 'mod', t.string_node(it.mod))
	to_object(obj, 'val', t.string_node(it.val))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	return obj
}

fn (t Tree) assoc(it ast.Assoc) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Assoc'))
	to_object(obj, 'var_name', t.string_node(it.var_name))
	s_arr := create_array()
	for f in it.fields {
		to_array(s_arr, t.string_node(f))
	}
	to_object(obj, 'fields', s_arr)
	e_arr := create_array()
	for e in it.exprs {
		to_array(e_arr, t.expr(e))
	}
	to_object(obj, 'exprs', e_arr)
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	return obj
}

fn (t Tree) cast_expr(it ast.CastExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('CastExpr'))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'arg', t.expr(it.arg))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'typname', t.string_node(it.typname))
	to_object(obj, 'expr_type', t.number_node(int(it.expr_type)))
	to_object(obj, 'has_arg', t.bool_node(it.has_arg))
	return obj
}

fn (t Tree) as_cast(it ast.AsCast) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('AsCast'))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'expr_type', t.number_node(int(it.expr_type)))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) type_expr(it ast.Type) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Type'))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	return obj
}

fn (t Tree) size_of(it ast.SizeOf) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('SizeOf'))
	to_object(obj, 'type_name', t.string_node(it.type_name))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	return obj
}

fn (t Tree) prefix_expr(it ast.PrefixExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('PrefixExpr'))
	to_object(obj, 'op', t.number_node(int(it.op)))
	to_object(obj, 'right', t.expr(it.right))
	return obj
}

fn (t Tree) assign_expr(it ast.AssignExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('AssignExpr'))
	to_object(obj, 'op', t.number_node(int(it.op)))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'left', t.expr(it.left))
	to_object(obj, 'val', t.expr(it.val))
	to_object(obj, 'left_type', t.number_node(int(it.left_type)))
	to_object(obj, 'right_type', t.number_node(int(it.right_type)))
	return obj
}

fn (t Tree) infix_expr(it ast.InfixExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('InfixExpr'))
	to_object(obj, 'op', t.number_node(int(it.op)))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'left', t.expr(it.left))
	to_object(obj, 'left_type', t.number_node(int(it.left_type)))
	to_object(obj, 'right', t.expr(it.right))
	to_object(obj, 'right_type', t.number_node(int(it.right_type)))
	return obj
}

fn (t Tree) index_expr(it ast.IndexExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('IndexExpr'))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'left', t.expr(it.left))
	to_object(obj, 'index', t.expr(it.index))
	to_object(obj, 'left_type', t.number_node(int(it.left_type)))
	to_object(obj, 'is_setter', t.bool_node(it.is_setter))
	return obj
}

fn (t Tree) postfix_expr(it ast.PostfixExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('PostfixExpr'))
	to_object(obj, 'op', t.number_node(int(it.op)))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) selector_expr(it ast.SelectorExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('SelectorExpr'))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'field_name', t.string_node(it.field_name))
	to_object(obj, 'expr_type', t.number_node(int(it.expr_type)))
	return obj
}

fn (t Tree) range_expr(it ast.RangeExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('RangeExpr'))
	to_object(obj, 'low', t.expr(it.low))
	to_object(obj, 'high', t.expr(it.high))
	return obj
}

fn (t Tree) if_expr(it ast.IfExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('IfExpr'))
	to_object(obj, 'tok_kind', t.number_node(int(it.tok_kind)))
	branch_arr := create_array()
	for b in it.branches {
		to_array(branch_arr, t.if_branch(b))
	}
	to_object(obj, 'branches', branch_arr)
	to_object(obj, 'left', t.expr(it.left))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'has_else', t.bool_node(it.has_else))
	to_object(obj, 'is_expr', t.bool_node(it.is_expr))
	return obj
}

fn (t Tree) if_branch(it ast.IfBranch) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('IfBranch'))
	to_object(obj, 'cond', t.expr(it.cond))
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'comment', t.comment(it.comment))
	return obj
}

fn (t Tree) ident(it ast.Ident) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Ident'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'value', t.string_node(it.value))
	to_object(obj, 'language', t.number_node(int(it.language)))
	to_object(obj, 'is_mut', t.bool_node(it.is_mut))
	to_object(obj, 'tok_kind', t.number_node(int(it.tok_kind)))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'kind', t.number_node(int(it.kind)))
	to_object(obj, 'info', t.ident_info(it.info))
	return obj
}

fn (t Tree) ident_info(info ast.IdentInfo) &C.cJSON {
	match info {
		ast.IdentVar { return t.ident_var(it) }
		ast.IdentFn { return t.ident_fn(it) }
	}
}

fn (t Tree) ident_var(it ast.IdentVar) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('IdentVar'))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'is_mut', t.bool_node(it.is_mut))
	to_object(obj, 'is_static', t.bool_node(it.is_static))
	to_object(obj, 'is_optional', t.bool_node(it.is_optional))
	return obj
}

fn (t Tree) ident_fn(it ast.IdentFn) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('IdentFn'))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	return obj
}

fn (t Tree) call_expr(it ast.CallExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('CallExpr'))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'left', t.expr(it.left))
	to_object(obj, 'is_method', t.bool_node(it.is_method))
	to_object(obj, 'mod', t.string_node(it.mod))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'language', t.number_node(int(it.language)))
	arg_arr := create_array()
	for e in it.args {
		to_array(arg_arr, t.call_arg(e))
	}
	to_object(obj, 'args', arg_arr)
	t_arr := create_array()
	for e in it.expected_arg_types {
		to_array(t_arr, t.number_node(int(e)))
	}
	to_object(obj, 'expected_arg_types', t_arr)
	to_object(obj, 'or_block', t.or_expr(it.or_block))
	to_object(obj, 'left_type', t.number_node(int(it.left_type)))
	to_object(obj, 'receiver_type', t.number_node(int(it.receiver_type)))
	to_object(obj, 'return_type', t.number_node(int(it.return_type)))
	to_object(obj, 'generic_type', t.number_node(int(it.generic_type)))
	return obj
}

fn (t Tree) call_arg(it ast.CallArg) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('CallArg'))
	to_object(obj, 'is_mut', t.bool_node(it.is_mut))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	return obj
}

fn (t Tree) or_expr(it ast.OrExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('OrExpr'))
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	to_object(obj, 'kind', t.number_node(int(it.kind)))
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) struct_init(it ast.StructInit) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('StructInit'))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'is_short', t.bool_node(it.is_short))
	s_arr := create_array()
	for f in it.fields {
		to_array(s_arr, t.struct_init_field(f))
	}
	to_object(obj, 'fields', s_arr)
	return obj
}

fn (t Tree) struct_init_field(it ast.StructInitField) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('StructInitField'))
	to_object(obj, 'name', t.string_node(it.name))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'expected_type', t.number_node(int(it.expected_type)))
	return obj
}

fn (t Tree) array_init(it ast.ArrayInit) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ArrayInit'))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	to_object(obj, 'elem_type', t.number_node(int(it.elem_type)))
	expr_arr := create_array()
	for e in it.exprs {
		to_array(expr_arr, t.expr(e))
	}
	to_object(obj, 'exprs', expr_arr)
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'elem_type_pos', t.position(it.elem_type_pos))
	to_object(obj, 'is_fixed', t.bool_node(it.is_fixed))
	to_object(obj, 'has_val', t.bool_node(it.has_val))
	to_object(obj, 'mod', t.string_node(it.mod))
	to_object(obj, 'len_expr', t.expr(it.len_expr))
	to_object(obj, 'cap_expr', t.expr(it.cap_expr))
	to_object(obj, 'default_expr', t.expr(it.default_expr))
	to_object(obj, 'has_len', t.bool_node(it.has_len))
	to_object(obj, 'has_cap', t.bool_node(it.has_cap))
	to_object(obj, 'has_default', t.bool_node(it.has_default))
	to_object(obj, 'is_interface', t.bool_node(it.is_interface))
	to_object(obj, 'interface_type', t.number_node(int(it.interface_type)))
	i_arr := create_array()
	for i in it.interface_types {
		to_array(i_arr, t.number_node(int(i)))
	}
	to_object(obj, 'interface_types', i_arr)
	return obj
}

fn (t Tree) map_init(it ast.MapInit) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('MapInit'))
	to_object(obj, 'typ', t.number_node(int(it.typ)))
	k_arr := create_array()
	for k in it.keys {
		to_array(k_arr, t.expr(k))
	}
	to_object(obj, 'keys', k_arr)
	v_arr := create_array()
	for v in it.vals {
		to_array(v_arr, t.expr(v))
	}
	to_object(obj, 'vals', v_arr)
	to_object(obj, 'pos', t.position(it.pos))
	return obj
}

fn (t Tree) none_expr(it ast.None) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('None'))
	// todo
	to_object(obj, 'foo', t.number_node(it.foo))
	return obj
}

fn (t Tree) par_expr(it ast.ParExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ParExpr'))
	to_object(obj, 'expr', t.expr(it.expr))
	return obj
}

fn (t Tree) if_guard_expr(it ast.IfGuardExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('IfGuardExpr'))
	to_object(obj, 'var_name', t.string_node(it.var_name))
	to_object(obj, 'expr', t.expr(it.expr))
	return obj
}

fn (t Tree) match_expr(it ast.MatchExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('MatchExpr'))
	to_object(obj, 'tok_kind', t.number_node(int(it.tok_kind)))
	to_object(obj, 'cond', t.expr(it.cond))
	m_arr := create_array()
	for b in it.branches {
		to_array(m_arr, t.match_branch(b))
	}
	to_object(obj, 'branches', m_arr)
	to_object(obj, 'cond_type', t.number_node(int(it.cond_type)))
	to_object(obj, 'return_type', t.number_node(int(it.return_type)))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'is_sum_type', t.bool_node(it.is_sum_type))
	to_object(obj, 'is_expr', t.bool_node(it.is_expr))
	to_object(obj, 'is_mut', t.bool_node(it.is_mut))
	return obj
}

fn (t Tree) match_branch(it ast.MatchBranch) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('MatchBranch'))
	expr_arr := create_array()
	for e in it.exprs {
		to_array(expr_arr, t.expr(e))
	}
	to_object(obj, 'exprs', expr_arr)
	stmt_arr := create_array()
	for s in it.stmts {
		to_array(stmt_arr, t.stmt(s))
	}
	to_object(obj, 'stmts', stmt_arr)
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'comment', t.comment(it.comment))
	to_object(obj, 'is_else', t.bool_node(it.is_else))
	return obj
}

fn (t Tree) concat_expr(it ast.ConcatExpr) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('ConcatExpr'))
	expr_arr := create_array()
	for e in it.vals {
		to_array(expr_arr, t.expr(e))
	}
	to_object(obj, 'vals', expr_arr)
	to_object(obj, 'return_type', t.number_node(int(it.return_type)))
	return obj
}

fn (t Tree) type_of(it ast.TypeOf) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('TypeOf'))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'expr_type', t.number_node(int(it.expr_type)))
	return obj
}

fn (t Tree) likely(it ast.Likely) &C.cJSON {
	obj := create_object()
	to_object(obj, 'ast_type', t.string_node('Likely'))
	to_object(obj, 'expr', t.expr(it.expr))
	to_object(obj, 'pos', t.position(it.pos))
	to_object(obj, 'is_likely', t.bool_node(it.is_likely))
	return obj
}

[inline]
fn to_object(node &C.cJSON, key string, child &C.cJSON) {
	add_item_to_object(node, key, child)
}

[inline]
fn to_array(node, child &C.cJSON) {
	add_item_to_array(node, child)
}

// get absolute path for file
fn abs_path(path string) string {
	if os.is_abs_path(path) {
		return path
	} else if path.starts_with('./') {
		return os.join_path(os.getwd(), path[2..])
	} else {
		return os.join_path(os.getwd(), path)
	}
}
